module Control(



);